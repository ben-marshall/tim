--! ------------------------------------------------------------------------------------------------
--!
--! @file tim_cpu_arch.vhdl
--! @brief Contains the architecture declaration/defintion for the TIM CPU module.
--!
--! ------------------------------------------------------------------------------------------------


--! Use the standard IEEE libraries
library ieee;
--! Import standard logic interfaces.
use ieee.std_logic_1164.ALL;
--! Standard numeric operations and types.
use ieee.numeric_std.ALL;
