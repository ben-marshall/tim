--! ------------------------------------------------------------------------------------------------
--!
--! @file bus_master.vhdl
--! @brief Source code for the master bus controller.
--!
--! ------------------------------------------------------------------------------------------------

