--! ------------------------------------------------------------------------------------------------
--!
--! @file top_synth.vhdl
--! @brief Top file for synthesised version of the TIM Processor.
--!
--! ------------------------------------------------------------------------------------------------
