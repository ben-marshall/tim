--! ------------------------------------------------------------------------------------------------
--!
--! @file mem_dummy.vhdl
--! @brief Source code for a dummy memory module used in simulations.
--!
--! ------------------------------------------------------------------------------------------------

