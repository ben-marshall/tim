--! ------------------------------------------------------------------------------------------------
--!
--! @file top_sim.vhdl
--! @brief Top file for simulated version of the TIM Processor.
--!
--! ------------------------------------------------------------------------------------------------
