--! ------------------------------------------------------------------------------------------------
--!
--! @file  bus_device_testbench.vhdl
--! @brief Contains the testbench for all bus devices.
--!
--! ------------------------------------------------------------------------------------------------

--! Use the standard IEEE libraries
library ieee;
--! Import standard logic interfaces.
use ieee.std_logic_1164.ALL;
--! Standard numeric operations and types.
use ieee.numeric_std.ALL;

