--! ------------------------------------------------------------------------------------------------
--!
--! @file alu.vhdl
--! @brief File containing source code for the basic ALU.
--!
--! ------------------------------------------------------------------------------------------------

