--! ------------------------------------------------------------------------------------------------
--!
--! @file sram_controller.vhdl
--! @brief Source code for the SRAM memory controller used in synthesis.
--!
--! ------------------------------------------------------------------------------------------------

