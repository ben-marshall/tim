--! ------------------------------------------------------------------------------------------------
--!
--! @file tim_cpu.vhdl
--! @brief Top file for the CPU module
--!
--! ------------------------------------------------------------------------------------------------

