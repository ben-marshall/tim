--! ------------------------------------------------------------------------------------------------
--!
--! @file bus_master_arch.vhdl
--! @brief Source code for the architecture declaration of the master bus controller.
--!
--! ------------------------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.ALL;
use ieee.numeric_std.ALL;

use work.tim_bus.tim_bus_data_width;
use work.tim_bus.tim_bus_burst_width;

architecture tim_bus_master_rtl of tim_bus_master is


begin


end architecture tim_bus_master_rtl;
