--! ------------------------------------------------------------------------------------------------
--!
--! @file  bus_device_master.vhdl
--! @brief Contains the architecture declaration of the master bus device. This architecture belongs
--!        to the bus_device entity.
--!
--! ------------------------------------------------------------------------------------------------

