--! ------------------------------------------------------------------------------------------------
--!
--! @file  bus_device_slave.vhdl
--! @brief Contains the architecture declaration of the slave bus device. This architecture belongs
--!        to the bus_device entity.
--!
--! ------------------------------------------------------------------------------------------------

