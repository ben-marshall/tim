--! ------------------------------------------------------------------------------------------------
--!
--! @file bus_slave.vhdl
--! @brief Source code for the slave bus controller.
--!
--! ------------------------------------------------------------------------------------------------

